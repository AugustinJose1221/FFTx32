`timescale 1ns/10ps
module FFTtb;

reg signed [11:0] r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31;
reg enable;
reg clk;
wire ret;
MyTestbed Test(.r0(r0),
	       .r1(r1),
	       .r2(r2),
	       .r3(r3),
	       .r4(r4),
	       .r5(r5),
	       .r6(r6),
	       .r7(r7),
	       .r8(r8),
	       .r9(r9),
	       .r10(r10),
	       .r11(r11),
	       .r12(r12),
	       .r13(r13),
	       .r14(r14),
	       .r15(r15),
	       .r16(r16),
	       .r17(r17),
	       .r18(r18),
	       .r19(r19),
	       .r20(r20),
	       .r21(r21),
	       .r22(r22),
	       .r23(r23),
	       .r24(r24),
	       .r25(r25),
	       .r26(r26),
	       .r27(r27),
	       .r28(r28),
	       .r29(r29),
	       .r30(r30),
	       .r31(r31),
	       .i0(i0),
	       .i1(i1),
	       .i2(i2),
	       .i3(i3),
	       .i4(i4),
	       .i5(i5),
	       .i6(i6),
	       .i7(i7),
	       .i8(i8),
	       .i9(i9),
	       .i10(i10),
	       .i11(i11),
	       .i12(i12),
	       .i13(i13),
	       .i14(i14),
	       .i15(i15),
	       .i16(i16),
	       .i17(i17),
	       .i18(i18),
	       .i19(i19),
	       .i20(i20),
	       .i21(i21),
	       .i22(i22),
	       .i23(i23),
	       .i24(i24),
	       .i25(i25),
	       .i26(i26),
	       .i27(i27),
	       .i28(i28),
	       .i29(i29),
	       .i30(i30),
	       .i31(i31),
	       .enable(enable),
	       .clk(clk),
	       .ret(ret));
	       
integer i;
parameter cycle = 10.0;
always #(cycle/2.0) clk = ~clk;
initial 
begin
	clk = 1;
	enable = 1;
	r0 = 0;
	r1 = -1700;
	r2 = -1605;
	r3 = 412;
	r4 = 1363;
	r5 = -115;
	r6 = -209;
	r7 = 277;
	r8 = 381;
	r9 = 736;
	r10 = -1086;
	r11 = 42;
	r12 = 1346;
	r13 = 1889;
	r14 = -978;
	r15 = 96;
	r16 = -227;
	r17 = -1409;
	r18 = 1979;
	r19 = -477;
	r20 = 299;
	r21 = -751;
	r22 = 1563;
	r23 = -968;
	r24 = -1552;
	r25 = -723;
	r26 = -484;
	r27 = -1781;
	r28 = 2043;
	r29 = -527;
	r30 = -701;
	r31 = 1502;

	i0 = -1884;
	i1 = 1674;
	i2 = 262;
	i3 = 1052;
	i4 = -6;
	i5 = 1818;
	i6 = -36;
	i7 = -1932;
	i8 = -203;
	i9 = -1591;
	i10 = -1760;
	i11 = 47;
	i12 = -1397;
	i13 = -145;
	i14 = -24;
	i15 = -743;
	i16 = 116;
	i17 = 1596;
	i18 = -98;
	i19 = -1501;
	i20 = 681;
	i21 = 1002;
	i22 = -1492;
	i23 = -1465;
	i24 = 121;
	i25 = 86;
	i26 = 393;
	i27 = -49;
	i28 = -1910;
	i29 = 621;
	i30 = 672;
	i31 = 2032;
end

always @(ret)
begin
	if(ret==1)begin
	enable = 0;
	#10;
	enable = 1;
	r0 = 1536;
	r1 = 592;
	r2 = -1210;
	r3 = 1962;
	r4 = -205;
	r5 = 638;
	r6 = -93;
	r7 = -475;
	r8 = 1753;
	r9 = -2022;
	r10 = 709;
	r11 = -752;
	r12 = -949;
	r13 = 1926;
	r14 = 1124;
	r15 = 592;
	r16 = 556;
	r17 = -1268;
	r18 = 1717;
	r19 = -12;
	r20 = -1852;
	r21 = 1560;
	r22 = 1590;
	r23 = 93;
	r24 = -955;
	r25 = -1710;
	r26 = 1889;
	r27 = -1212;
	r28 = -286;
	r29 = 912;
	r30 = 1079;
	r31 = -605;

	i0 = -1427;
	i1 = -973;
	i2 = 1864;
	i3 = 1620;
	i4 = 488;
	i5 = -1410;
	i6 = 1042;
	i7 = 1644;
	i8 = -1037;
	i9 = 1093;
	i10 = 865;
	i11 = 46;
	i12 = 1805;
	i13 = -1718;
	i14 = 1519;
	i15 = 1587;
	i16 = 1748;
	i17 = -1915;
	i18 = -1195;
	i19 = -1887;
	i20 = -1765;
	i21 = 553;
	i22 = 970;
	i23 = 1382;
	i24 = -167;
	i25 = -1769;
	i26 = -950;
	i27 = -1066;
	i28 = -1922;
	i29 = -1630;
	i30 = -1256;
	i31 = -608;	
	end	
end

initial
begin
	$dumpfile("main.vcd");
	$dumpvars(0, FFTtb);
	#2050;
	$finish;
	
end



endmodule
					
		

	
